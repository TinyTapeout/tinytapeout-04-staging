VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_loopback
  CLASS BLOCK ;
  FOREIGN tt_um_loopback ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.550 2.480 44.150 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.145 2.480 84.745 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.740 2.480 125.340 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.335 2.480 165.935 106.320 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.255 2.480 23.855 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.850 2.480 64.450 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.445 2.480 105.045 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.040 2.480 145.640 106.320 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 107.800 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 107.800 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 107.260 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 107.800 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 107.800 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 107.800 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 107.260 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 107.260 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 105.900 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 107.260 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 107.800 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 107.800 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 107.800 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 107.800 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 107.800 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 107.800 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 107.800 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 107.800 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 105.220 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 103.180 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 105.220 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 107.260 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 105.220 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 105.220 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 105.220 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 105.220 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 107.260 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 105.220 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 105.220 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 105.220 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 105.900 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 105.220 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 105.220 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 105.220 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 105.900 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 105.900 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 107.260 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 103.180 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 105.900 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 105.900 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 103.180 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 107.260 66.850 108.800 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 101.945 165.330 104.775 ;
        RECT 2.570 96.505 165.330 99.335 ;
        RECT 2.570 91.065 165.330 93.895 ;
        RECT 2.570 85.625 165.330 88.455 ;
        RECT 2.570 80.185 165.330 83.015 ;
        RECT 2.570 74.745 165.330 77.575 ;
        RECT 2.570 69.305 165.330 72.135 ;
        RECT 2.570 63.865 165.330 66.695 ;
        RECT 2.570 58.425 165.330 61.255 ;
        RECT 2.570 52.985 165.330 55.815 ;
        RECT 2.570 47.545 165.330 50.375 ;
        RECT 2.570 42.105 165.330 44.935 ;
        RECT 2.570 36.665 165.330 39.495 ;
        RECT 2.570 31.225 165.330 34.055 ;
        RECT 2.570 25.785 165.330 28.615 ;
        RECT 2.570 20.345 165.330 23.175 ;
        RECT 2.570 14.905 165.330 17.735 ;
        RECT 2.570 9.465 165.330 12.295 ;
        RECT 2.570 4.025 165.330 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 165.140 106.165 ;
      LAYER met1 ;
        RECT 2.760 2.480 165.935 108.760 ;
      LAYER met2 ;
        RECT 7.910 2.535 165.905 108.790 ;
      LAYER met3 ;
        RECT 7.630 2.555 165.925 107.265 ;
      LAYER met4 ;
        RECT 8.370 104.820 10.950 107.265 ;
        RECT 12.050 104.820 14.630 107.265 ;
        RECT 15.730 104.820 18.310 107.265 ;
        RECT 19.410 106.860 21.990 107.265 ;
        RECT 23.090 106.860 25.670 107.265 ;
        RECT 19.410 106.720 25.670 106.860 ;
        RECT 19.410 104.820 21.855 106.720 ;
        RECT 7.655 102.855 21.855 104.820 ;
        RECT 24.255 104.820 25.670 106.720 ;
        RECT 26.770 104.820 29.350 107.265 ;
        RECT 24.255 102.855 29.350 104.820 ;
        RECT 30.450 104.820 33.030 107.265 ;
        RECT 34.130 104.820 36.710 107.265 ;
        RECT 37.810 104.820 40.390 107.265 ;
        RECT 41.490 106.720 44.070 107.265 ;
        RECT 41.490 104.820 42.150 106.720 ;
        RECT 45.170 105.500 47.750 107.265 ;
        RECT 48.850 105.500 51.430 107.265 ;
        RECT 45.170 104.820 51.430 105.500 ;
        RECT 52.530 104.820 55.110 107.265 ;
        RECT 56.210 104.820 58.790 107.265 ;
        RECT 59.890 106.860 62.470 107.265 ;
        RECT 63.570 106.860 66.150 107.265 ;
        RECT 67.250 106.860 69.830 107.265 ;
        RECT 59.890 106.720 69.830 106.860 ;
        RECT 59.890 104.820 62.450 106.720 ;
        RECT 30.450 102.855 42.150 104.820 ;
        RECT 44.550 102.855 62.450 104.820 ;
        RECT 64.850 102.855 69.830 106.720 ;
        RECT 70.930 105.500 73.510 107.265 ;
        RECT 74.610 105.500 77.190 107.265 ;
        RECT 78.290 105.500 80.870 107.265 ;
        RECT 70.930 102.855 80.870 105.500 ;
        RECT 81.970 106.860 84.550 107.265 ;
        RECT 85.650 106.860 88.230 107.265 ;
        RECT 81.970 106.720 88.230 106.860 ;
        RECT 81.970 102.855 82.745 106.720 ;
        RECT 85.145 105.500 88.230 106.720 ;
        RECT 89.330 105.500 91.910 107.265 ;
        RECT 93.010 106.860 125.030 107.265 ;
        RECT 126.130 106.860 128.710 107.265 ;
        RECT 93.010 106.720 128.710 106.860 ;
        RECT 93.010 105.500 103.045 106.720 ;
        RECT 85.145 102.855 103.045 105.500 ;
        RECT 105.445 102.855 123.340 106.720 ;
        RECT 125.740 105.500 128.710 106.720 ;
        RECT 129.810 106.860 132.390 107.265 ;
        RECT 133.490 106.860 136.070 107.265 ;
        RECT 137.170 106.860 150.790 107.265 ;
        RECT 129.810 106.720 151.505 106.860 ;
        RECT 129.810 105.500 143.640 106.720 ;
        RECT 125.740 102.855 143.640 105.500 ;
        RECT 146.040 102.855 151.505 106.720 ;
  END
END tt_um_loopback
END LIBRARY

