VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_marno_factorize
  CLASS BLOCK ;
  FOREIGN tt_um_marno_factorize ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.550 2.480 44.150 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.145 2.480 84.745 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.740 2.480 125.340 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.335 2.480 165.935 106.320 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.255 2.480 23.855 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.850 2.480 64.450 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.445 2.480 105.045 106.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.040 2.480 145.640 106.320 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 106.950 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 107.260 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 107.260 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 107.260 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 107.260 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 107.260 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 107.260 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 107.260 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 107.260 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 107.260 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 107.800 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 107.800 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 107.800 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 107.800 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 107.800 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 107.800 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 107.800 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 107.800 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 105.900 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 107.260 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 105.900 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 107.260 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 107.260 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 107.260 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 107.260 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 107.260 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 107.260 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 105.900 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 107.260 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 105.900 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 107.260 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 107.260 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 107.260 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 105.900 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 107.260 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 106.580 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 107.260 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 107.260 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 107.260 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 106.580 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 107.260 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 105.220 66.850 108.800 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 101.945 165.330 104.775 ;
        RECT 2.570 96.505 165.330 99.335 ;
        RECT 2.570 91.065 165.330 93.895 ;
        RECT 2.570 85.625 165.330 88.455 ;
        RECT 2.570 80.185 165.330 83.015 ;
        RECT 2.570 74.745 165.330 77.575 ;
        RECT 2.570 69.305 165.330 72.135 ;
        RECT 2.570 63.865 165.330 66.695 ;
        RECT 2.570 58.425 165.330 61.255 ;
        RECT 2.570 52.985 165.330 55.815 ;
        RECT 2.570 47.545 165.330 50.375 ;
        RECT 2.570 42.105 165.330 44.935 ;
        RECT 2.570 36.665 165.330 39.495 ;
        RECT 2.570 31.225 165.330 34.055 ;
        RECT 2.570 25.785 165.330 28.615 ;
        RECT 2.570 20.345 165.330 23.175 ;
        RECT 2.570 14.905 165.330 17.735 ;
        RECT 2.570 9.465 165.330 12.295 ;
        RECT 2.570 4.025 165.330 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 165.140 106.165 ;
      LAYER met1 ;
        RECT 2.760 2.480 165.935 107.400 ;
      LAYER met2 ;
        RECT 5.610 2.535 165.905 107.430 ;
      LAYER met3 ;
        RECT 5.585 2.555 165.925 107.265 ;
      LAYER met4 ;
        RECT 8.370 106.860 10.950 107.265 ;
        RECT 12.050 106.860 14.630 107.265 ;
        RECT 15.730 106.860 18.310 107.265 ;
        RECT 19.410 106.860 21.990 107.265 ;
        RECT 23.090 106.860 25.670 107.265 ;
        RECT 7.655 106.720 25.670 106.860 ;
        RECT 7.655 89.255 21.855 106.720 ;
        RECT 24.255 105.500 25.670 106.720 ;
        RECT 26.770 106.860 29.350 107.265 ;
        RECT 30.450 106.860 33.030 107.265 ;
        RECT 26.770 105.500 33.030 106.860 ;
        RECT 34.130 105.500 36.710 107.265 ;
        RECT 37.810 106.860 40.390 107.265 ;
        RECT 41.490 106.860 44.070 107.265 ;
        RECT 45.170 106.860 47.750 107.265 ;
        RECT 48.850 106.860 51.430 107.265 ;
        RECT 37.810 106.720 51.430 106.860 ;
        RECT 37.810 105.500 42.150 106.720 ;
        RECT 24.255 89.255 42.150 105.500 ;
        RECT 44.550 105.500 51.430 106.720 ;
        RECT 52.530 106.860 55.110 107.265 ;
        RECT 56.210 106.860 58.790 107.265 ;
        RECT 52.530 105.500 58.790 106.860 ;
        RECT 59.890 106.860 62.470 107.265 ;
        RECT 63.570 106.860 66.150 107.265 ;
        RECT 59.890 106.720 66.150 106.860 ;
        RECT 59.890 105.500 62.450 106.720 ;
        RECT 44.550 89.255 62.450 105.500 ;
        RECT 64.850 104.820 66.150 106.720 ;
        RECT 67.250 106.860 69.830 107.265 ;
        RECT 70.930 106.860 73.510 107.265 ;
        RECT 67.250 106.180 73.510 106.860 ;
        RECT 74.610 106.860 77.190 107.265 ;
        RECT 78.290 106.860 80.870 107.265 ;
        RECT 81.970 106.860 84.550 107.265 ;
        RECT 85.650 106.860 88.230 107.265 ;
        RECT 74.610 106.720 88.230 106.860 ;
        RECT 74.610 106.180 82.745 106.720 ;
        RECT 67.250 104.820 82.745 106.180 ;
        RECT 64.850 89.255 82.745 104.820 ;
        RECT 85.145 106.180 88.230 106.720 ;
        RECT 89.330 106.860 91.910 107.265 ;
        RECT 93.010 106.860 125.030 107.265 ;
        RECT 126.130 106.860 128.710 107.265 ;
        RECT 129.810 106.860 132.390 107.265 ;
        RECT 133.490 106.860 136.070 107.265 ;
        RECT 137.170 106.860 139.750 107.265 ;
        RECT 140.850 106.860 143.430 107.265 ;
        RECT 144.530 106.860 147.110 107.265 ;
        RECT 148.210 106.860 150.790 107.265 ;
        RECT 151.890 106.860 154.470 107.265 ;
        RECT 155.570 106.860 158.150 107.265 ;
        RECT 89.330 106.720 158.150 106.860 ;
        RECT 89.330 106.180 103.045 106.720 ;
        RECT 85.145 89.255 103.045 106.180 ;
        RECT 105.445 89.255 123.340 106.720 ;
        RECT 125.740 89.255 143.640 106.720 ;
        RECT 146.040 106.550 158.150 106.720 ;
        RECT 146.040 89.255 158.865 106.550 ;
  END
END tt_um_marno_factorize
END LIBRARY

